netcdf pf_active_coil_current {

// Global attributes
:title = "PF Active Coil Current" ;
:institution = "ITER Organization" ;
:source = "IMAS pf_active IDS current subset" ;
:conventions = "CF-1.8, IMAS-3.0" ;
:comment = "Poloidal field coil current time series and control data" ;

dimensions:
    // Time series dimensions
    time = _ ;                      // Number of time points
    coil = _ ;                      // Number of PF coils
    // Circuit topology dimensions
    circuit = _ ;                   // Number of independent circuits
    circuit_coil = _ ;              // Circuit-coil connections

variables:
    // Time coordinate
    double time(time) ;
        time:units = "s" ;
        time:long_name = "time coordinate" ;
        time:standard_name = "time" ;
        time:axis = "T" ;
        time:_FillValue = _ ;
        
    // Coil identifiers
    string coil_name(coil) ;
        coil_name:long_name = "coil identifier name" ;
        coil_name:description = "Human readable coil identifier (e.g., PF1, PF2, etc.)" ;

    // Circuit identifiers  
    string circuit_name(circuit) ;
        circuit_name:long_name = "circuit identifier name" ;
        circuit_name:description = "Power supply circuit identifier" ;

    // Current data
    double coil_current(time, coil) ;
        coil_current:units = "A" ;
        coil_current:long_name = "PF coil current" ;
        coil_current:standard_name = "electric_current" ;
        coil_current:coordinates = "time" ;
        coil_current:_FillValue = _ ;
        coil_current:description = "Time-dependent current in each PF coil" ;

    double circuit_current(time, circuit) ;
        circuit_current:units = "A" ;
        circuit_current:long_name = "PF circuit current" ;
        circuit_current:standard_name = "electric_current" ;
        circuit_current:coordinates = "time" ;
        circuit_current:_FillValue = _ ;
        circuit_current:description = "Time-dependent current in each independent circuit" ;

    // Circuit topology mapping
    int circuit_coil_index(circuit_coil) ;
        circuit_coil_index:long_name = "coil index for circuit connection" ;
        circuit_coil_index:description = "Maps circuit elements to coil indices" ;
        circuit_coil_index:valid_range = _, _ ;

    int circuit_index(circuit_coil) ;
        circuit_index:long_name = "circuit index for circuit connection" ;
        circuit_index:description = "Maps circuit elements to circuit indices" ;
        circuit_index:valid_range = _, _ ;

    double circuit_coil_turns(circuit_coil) ;
        circuit_coil_turns:units = "1" ;
        circuit_coil_turns:long_name = "number of turns in circuit-coil connection" ;
        circuit_coil_turns:description = "Turn ratio between circuit and coil" ;
        circuit_coil_turns:valid_min = _ ;

    // Control and reference data
    double coil_current_reference(time, coil) ;
        coil_current_reference:units = "A" ;
        coil_current_reference:long_name = "PF coil reference current" ;
        coil_current_reference:standard_name = "electric_current" ;
        coil_current_reference:coordinates = "time" ;
        coil_current_reference:_FillValue = _ ;
        coil_current_reference:description = "Commanded/reference current for PF coils" ;

    double circuit_voltage(time, circuit) ;
        circuit_voltage:units = "V" ;
        circuit_voltage:long_name = "PF circuit voltage" ;
        circuit_voltage:standard_name = "electric_potential_difference" ;
        circuit_voltage:coordinates = "time" ;
        circuit_voltage:_FillValue = _ ;
        circuit_voltage:description = "Time-dependent voltage across each circuit" ;

    // Electrical properties
    double coil_resistance(coil) ;
        coil_resistance:units = "Ohm" ;
        coil_resistance:long_name = "PF coil resistance" ;
        coil_resistance:description = "DC resistance of each coil" ;
        coil_resistance:valid_min = _ ;

    double coil_inductance(coil) ;
        coil_inductance:units = "H" ;
        coil_inductance:long_name = "PF coil self-inductance" ;
        coil_inductance:description = "Self-inductance of each coil" ;
        coil_inductance:valid_min = _ ;

    // Power and energy
    double coil_power(time, coil) ;
        coil_power:units = "W" ;
        coil_power:long_name = "PF coil power consumption" ;
        coil_power:coordinates = "time" ;
        coil_power:_FillValue = _ ;
        coil_power:description = "Instantaneous power consumption in each coil" ;

    double circuit_energy(time, circuit) ;
        circuit_energy:units = "J" ;
        circuit_energy:long_name = "PF circuit stored energy" ;
        circuit_energy:coordinates = "time" ;
        circuit_energy:_FillValue = _ ;
        circuit_energy:description = "Magnetic energy stored in each circuit" ;
}
