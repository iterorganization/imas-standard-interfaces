netcdf tf_active_coil_geometry {

// Global attributes
:title = "TF Active Coil Geometry" ;
:institution = "ITER Organization" ;
:source = "IMAS tf_active IDS geometry subset" ;
:conventions = "CF-1.8, IMAS-3.0" ;
:comment = "Toroidal field coil geometric description including 3D geometry containers" ;

dimensions:
    // Coil structure dimensions
    coil = UNLIMITED ;                      // Number of TF coils (typically 18 for ITER)
    toroidal_angle = UNLIMITED ;            // Number of toroidal positions
      // TF outline geometry dimensions (poloidal cross-section)
    tf_outline_node = UNLIMITED ;           // Nodes for coil outlines  
    tf_outline_element = UNLIMITED ;        // Number of outline elements (one per coil)
    
    // TF 3D element geometry dimensions
    tf_element_node = UNLIMITED ;           // Nodes for 3D coil elements
    tf_element = UNLIMITED ;                // Total number of 3D coil elements

variables:    // Toroidal angle coordinate
    double toroidal_angle(toroidal_angle) ;
        toroidal_angle:units = "rad" ;
        toroidal_angle:long_name = "toroidal angle coordinate" ;
        toroidal_angle:standard_name = "angle" ;
        toroidal_angle:axis = "Z" ;

    // Coil identifiers
    string coil_name(coil) ;
        coil_name:long_name = "coil identifier name" ;
        coil_name:description = "Human readable coil identifier (e.g., TF01, TF02, etc.)" ;

    // TF outline geometry container (2D poloidal cross-section)
    int tf_outline_geometry ;
        tf_outline_geometry:geometry_type = "polygon" ;
        tf_outline_geometry:node_coordinates = "tf_outline_r tf_outline_z" ;
        tf_outline_geometry:node_count = "tf_outline_node_count" ;
        tf_outline_geometry:coordinates = "tf_outline_r tf_outline_z" ;
        tf_outline_geometry:description = "TF coil outline geometry container (poloidal cross-section)" ;    // TF outline coordinate variables
    double tf_outline_r(tf_outline_node) ;
        tf_outline_r:units = "m" ;
        tf_outline_r:long_name = "TF outline major radius coordinate" ;
        tf_outline_r:standard_name = "projection_r_coordinate" ;

    double tf_outline_z(tf_outline_node) ;
        tf_outline_z:units = "m" ;
        tf_outline_z:long_name = "TF outline vertical coordinate" ;
        tf_outline_z:standard_name = "projection_z_coordinate" ;

    // TF outline topology
    int tf_outline_node_count(tf_outline_element) ;
        tf_outline_node_count:long_name = "number of nodes per TF outline element" ;
        tf_outline_node_count:description = "Node count for each coil outline polygon" ;    int tf_outline_coil_index(tf_outline_element) ;
        tf_outline_coil_index:long_name = "coil index for TF outline element" ;
        tf_outline_coil_index:description = "Maps outline elements to parent coil" ;
        tf_outline_coil_index:valid_min = 0 ;

    // TF 3D element geometry container
    int tf_element_geometry ;
        tf_element_geometry:geometry_type = "polygon" ;
        tf_element_geometry:node_coordinates = "tf_element_r tf_element_z tf_element_phi" ;
        tf_element_geometry:node_count = "tf_element_node_count" ;
        tf_element_geometry:coordinates = "tf_element_r tf_element_z tf_element_phi" ;
        tf_element_geometry:description = "3D TF coil element geometry container" ;    // TF 3D element coordinate variables
    double tf_element_r(tf_element_node) ;
        tf_element_r:units = "m" ;
        tf_element_r:long_name = "TF element major radius coordinate" ;
        tf_element_r:standard_name = "projection_r_coordinate" ;

    double tf_element_z(tf_element_node) ;
        tf_element_z:units = "m" ;
        tf_element_z:long_name = "TF element vertical coordinate" ;
        tf_element_z:standard_name = "projection_z_coordinate" ;

    double tf_element_phi(tf_element_node) ;
        tf_element_phi:units = "rad" ;
        tf_element_phi:long_name = "TF element toroidal angle coordinate" ;
        tf_element_phi:standard_name = "angle" ;

    // TF 3D element topology
    int tf_element_node_count(tf_element) ;
        tf_element_node_count:long_name = "number of nodes per TF 3D element" ;
        tf_element_node_count:description = "Node count for each 3D element polygon" ;    int tf_element_coil_index(tf_element) ;
        tf_element_coil_index:long_name = "coil index for TF element" ;
        tf_element_coil_index:description = "Maps 3D elements to parent coil" ;
        tf_element_coil_index:valid_min = 0 ;

    int tf_element_poloidal_index(tf_element) ;
        tf_element_poloidal_index:long_name = "poloidal segment index for TF element" ;
        tf_element_poloidal_index:description = "Poloidal subdivision index within coil" ;
        tf_element_poloidal_index:valid_min = 0 ;

    int tf_element_toroidal_index(tf_element) ;
        tf_element_toroidal_index:long_name = "toroidal segment index for TF element" ;
        tf_element_toroidal_index:description = "Toroidal subdivision index within coil" ;
        tf_element_toroidal_index:valid_min = 0 ;

    // Geometric properties
    double coil_volume(coil) ;
        coil_volume:units = "m^3" ;
        coil_volume:long_name = "total coil volume" ;
        coil_volume:description = "Sum of all 3D element volumes for each coil" ;

    double tf_element_volume(tf_element) ;
        tf_element_volume:units = "m^3" ;
        tf_element_volume:long_name = "TF element volume" ;
        tf_element_volume:geometry = "tf_element_geometry" ;

    // Coil center coordinates
    double coil_center_r(coil) ;
        coil_center_r:units = "m" ;
        coil_center_r:long_name = "coil geometric center major radius" ;
        coil_center_r:description = "Volume-weighted center of coil elements" ;

    double coil_center_z(coil) ;
        coil_center_z:units = "m" ;
        coil_center_z:long_name = "coil geometric center vertical coordinate" ;
        coil_center_z:description = "Volume-weighted center of coil elements" ;

    double coil_center_phi(coil) ;
        coil_center_phi:units = "rad" ;
        coil_center_phi:long_name = "coil geometric center toroidal angle" ;
        coil_center_phi:description = "Volume-weighted center toroidal position" ;    // Magnetic properties  
    double coil_turns(coil) ;
        coil_turns:units = "1" ;
        coil_turns:long_name = "number of turns per TF coil" ;
        coil_turns:description = "Total number of conductor turns in each coil" ;
        coil_turns:valid_min = 0.0 ;

    double coil_current_density(coil) ;
        coil_current_density:units = "A/m^2" ;
        coil_current_density:long_name = "coil current density" ;
        coil_current_density:description = "Average current density in coil conductor" ;
}
